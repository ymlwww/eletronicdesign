library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity plant is
	port(
		 plantkind: in std_logic_vector(4 downto 0);
		 lifetime: out std_logic_vector(6 downto 0);
		 recovertime: out std_logic_vector(5 downto 0);
		 fire: out std_logic_vector(6 downto 0);
		 fireinterval: out std_logic_vector(3 downto 0);
		 fireradius: out std_logic_vector(6 downto 0);
		 price: out std_logic_vector(6 downto 0);
		 sunariseinterval: out std_logic_vector(5 downto 0);
		 preparetime: out std_logic_vector(5 downto 0);
		 address:out std_logic_vector(18 downto 0); --注意加零
		 --address的具体每位分布待定
		 lasttime:out std_logic_vector(3 downto 0)
	);
end plant;

architecture plantbehavioral of plant is
	signal addressinfo:std_logic_vector(31 downto 0);
	--address info：前一位存储植物的生命值，生命值一般植物生命值3，南瓜和坚果80；
	--第二位到第四位存储植物的价格，价格有25,50,100,125,150,175,一共六种
	--第五位存储植物的攻击力，一共两种，20,1800；
	--第六位存储冷却时间，一共两种，8,30，50改三十；
	--第七位到第九位存储时间间隔，有2（攻击间隔）,24(阳光产生间隔),4,15,42,1,一共六种
	--第十一位到第十三位存储攻击范围，有前方一整行，2格半径，单行前后两格，正前方2格，前后2格，三整行，前后一个，一整行，一共六种
	--剩下十九位存储动画的的开头地址，默认每个动画是5帧，也就是一共是5个连续的地址
begin	
	--读取sram
	--process(address) --此部分内容有待sram读写程序完善
	--此process的目的在于读取sram
	--begin
	--此部分需要对addressinfo赋值
	--end process;
	process(plantkind,address,addressinfo)
	--首先是根据plantkind得出对应的address的位置
	--其次是根据address读出adressinfo
	if(addressinfo[0] = '1')
		lifetime<="1010000";
	else
		lifetime<="0000011";
	case addressinfo(1 to 3) is
		when 
	
	
end plantbehavioral;
